`timescale 1ns / 100ps
`define SEED    'h1AA

module tb_filter();

    parameter SEED = `SEED;

    reg clock;
    reg i_reset;
    wire reset;

    
    wire                  valid                   ;
    wire                  prbs9_out               ;
    wire signed [7:0]     filter_out              ;

    reg  signed [7:0]     rx_buffer        [3:0]  ;
    wire                  rx_bit                  ; 

    wire signed [0:7]     expected_output  [0:799];
    wire signed [0:7]     expected_sample         ;
    wire                  expected_bit            ;
    wire        [0:799]   expected_rx_bits = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b0,1'b0};
    
    reg   [10:0]          ptr1                    ;
    reg   [10:0]          ptr2                    ;
    reg   [10:0]          ptr3                    ;

    reg   [63:0]          error_count_samples     ; //! error count for samples
    reg   [63:0]          error_count             ; //! error count
    

    initial
    begin
        clock               = 1'b0       ;  // inicializo clock
        i_reset             = 1'b0       ;  // activo reset (activo por bajo)
        
        // en t = 100 ns
        #100 i_reset        = 1'b1       ;  // desactivo el reset
    end

    always #5 clock = ~clock; // 5ns en bajo y 5ns en alto, periodo de 10ns

    integer i;
    always @(posedge clock) 
        begin
            if (reset)
                begin
                    error_count <= 0;
                    error_count_samples <= 0;
                    ptr1 <= 0;
                    ptr2 <= 0;
                    ptr3 <= 0;
                end
            else
                begin                    
                    // shift buffer de entrada
                    rx_buffer[0] <= filter_out;

                    for (i = 1; i < 4; i=i+1)
                        rx_buffer[i] <= rx_buffer[i-1];
                 
                        
                    // comparo con valores esperados
                    ptr3 <= ptr3 + 1;
                    
                    if (ptr3 > 3) // delay
                    begin
                        ptr2 <= ptr2 + 1;
                        if (filter_out != expected_sample)
                            error_count_samples <= error_count_samples + 1;
                    end

                    if (ptr3 > 4) // delay, una mas por el buffer_rx
                    begin
                        ptr1 <= ptr1 + 1;
                        if (rx_bit != expected_bit)
                            error_count <= error_count + 1;
                    end

                    if (ptr2 == 800)
                    begin
                        $display("Error count bits: %d", error_count);
                        $display("Error count samples %d", error_count_samples);
                        $finish;
                    end
                end
        end
    
    prbs9 # (
        .SEED   (SEED)
    )
        u_prbs9 (
            .o_bit      (prbs9_out)     ,
            .i_enable   (valid)         ,
            .i_reset    (reset)         ,
            .clock      (clock)     
        );

    control #(
            .NB_COUNT (2)
        )
        u_control (
            .o_valid  (valid)     ,
            .i_reset  (reset)     ,
            .clock    (clock)
        );

    filter #()
        u_filter (
            .i_enable  (i_reset)   ,
            .i_valid   (valid)     ,
            .i_bit     (prbs9_out) ,
            .o_data     (filter_out),
            .reset     (reset)     ,
            .clock     (clock)
        );

    
    assign rx_bit = rx_buffer[0][7];
    assign expected_bit     = expected_rx_bits[ptr1];
    assign expected_sample  = expected_output[ptr2];
    assign reset    = ~i_reset        ;


    assign expected_output[0] = 8'd126;
    assign expected_output[1] = 8'd124;
    assign expected_output[2] = 8'd120;
    assign expected_output[3] = 8'd120;
    assign expected_output[4] = 8'd124;
    assign expected_output[5] = 8'd127;
    assign expected_output[6] = 8'd127;
    assign expected_output[7] = 8'd127;
    assign expected_output[8] = 8'd127;
    assign expected_output[9] = 8'd58;
    assign expected_output[10] = 8'd224;
    assign expected_output[11] = 8'd150;
    assign expected_output[12] = 8'd128;
    assign expected_output[13] = 8'd170;
    assign expected_output[14] = 8'd4;
    assign expected_output[15] = 8'd90;
    assign expected_output[16] = 8'd127;
    assign expected_output[17] = 8'd90;
    assign expected_output[18] = 8'd0;
    assign expected_output[19] = 8'd166;
    assign expected_output[20] = 8'd128;
    assign expected_output[21] = 8'd166;
    assign expected_output[22] = 8'd0;
    assign expected_output[23] = 8'd90;
    assign expected_output[24] = 8'd127;
    assign expected_output[25] = 8'd90;
    assign expected_output[26] = 8'd0;
    assign expected_output[27] = 8'd166;
    assign expected_output[28] = 8'd130;
    assign expected_output[29] = 8'd166;
    assign expected_output[30] = 8'd252;
    assign expected_output[31] = 8'd86;
    assign expected_output[32] = 8'd126;
    assign expected_output[33] = 8'd106;
    assign expected_output[34] = 8'd36;
    assign expected_output[35] = 8'd202;
    assign expected_output[36] = 8'd130;
    assign expected_output[37] = 8'd128;
    assign expected_output[38] = 8'd128;
    assign expected_output[39] = 8'd128;
    assign expected_output[40] = 8'd128;
    assign expected_output[41] = 8'd186;
    assign expected_output[42] = 8'd4;
    assign expected_output[43] = 8'd74;
    assign expected_output[44] = 8'd126;
    assign expected_output[45] = 8'd127;
    assign expected_output[46] = 8'd127;
    assign expected_output[47] = 8'd127;
    assign expected_output[48] = 8'd127;
    assign expected_output[49] = 8'd120;
    assign expected_output[50] = 8'd116;
    assign expected_output[51] = 8'd120;
    assign expected_output[52] = 8'd126;
    assign expected_output[53] = 8'd127;
    assign expected_output[54] = 8'd127;
    assign expected_output[55] = 8'd127;
    assign expected_output[56] = 8'd126;
    assign expected_output[57] = 8'd74;
    assign expected_output[58] = 8'd4;
    assign expected_output[59] = 8'd186;
    assign expected_output[60] = 8'd130;
    assign expected_output[61] = 8'd128;
    assign expected_output[62] = 8'd128;
    assign expected_output[63] = 8'd128;
    assign expected_output[64] = 8'd128;
    assign expected_output[65] = 8'd202;
    assign expected_output[66] = 8'd32;
    assign expected_output[67] = 8'd102;
    assign expected_output[68] = 8'd127;
    assign expected_output[69] = 8'd102;
    assign expected_output[70] = 8'd28;
    assign expected_output[71] = 8'd198;
    assign expected_output[72] = 8'd132;
    assign expected_output[73] = 8'd128;
    assign expected_output[74] = 8'd128;
    assign expected_output[75] = 8'd128;
    assign expected_output[76] = 8'd128;
    assign expected_output[77] = 8'd136;
    assign expected_output[78] = 8'd140;
    assign expected_output[79] = 8'd136;
    assign expected_output[80] = 8'd132;
    assign expected_output[81] = 8'd128;
    assign expected_output[82] = 8'd128;
    assign expected_output[83] = 8'd128;
    assign expected_output[84] = 8'd128;
    assign expected_output[85] = 8'd198;
    assign expected_output[86] = 8'd32;
    assign expected_output[87] = 8'd106;
    assign expected_output[88] = 8'd127;
    assign expected_output[89] = 8'd86;
    assign expected_output[90] = 8'd0;
    assign expected_output[91] = 8'd170;
    assign expected_output[92] = 8'd130;
    assign expected_output[93] = 8'd150;
    assign expected_output[94] = 8'd220;
    assign expected_output[95] = 8'd54;
    assign expected_output[96] = 8'd126;
    assign expected_output[97] = 8'd127;
    assign expected_output[98] = 8'd127;
    assign expected_output[99] = 8'd127;
    assign expected_output[100] = 8'd127;
    assign expected_output[101] = 8'd70;
    assign expected_output[102] = 8'd0;
    assign expected_output[103] = 8'd186;
    assign expected_output[104] = 8'd130;
    assign expected_output[105] = 8'd128;
    assign expected_output[106] = 8'd128;
    assign expected_output[107] = 8'd128;
    assign expected_output[108] = 8'd128;
    assign expected_output[109] = 8'd202;
    assign expected_output[110] = 8'd32;
    assign expected_output[111] = 8'd102;
    assign expected_output[112] = 8'd127;
    assign expected_output[113] = 8'd102;
    assign expected_output[114] = 8'd28;
    assign expected_output[115] = 8'd198;
    assign expected_output[116] = 8'd130;
    assign expected_output[117] = 8'd128;
    assign expected_output[118] = 8'd128;
    assign expected_output[119] = 8'd128;
    assign expected_output[120] = 8'd128;
    assign expected_output[121] = 8'd128;
    assign expected_output[122] = 8'd128;
    assign expected_output[123] = 8'd128;
    assign expected_output[124] = 8'd130;
    assign expected_output[125] = 8'd182;
    assign expected_output[126] = 8'd252;
    assign expected_output[127] = 8'd70;
    assign expected_output[128] = 8'd126;
    assign expected_output[129] = 8'd127;
    assign expected_output[130] = 8'd127;
    assign expected_output[131] = 8'd127;
    assign expected_output[132] = 8'd127;
    assign expected_output[133] = 8'd54;
    assign expected_output[134] = 8'd224;
    assign expected_output[135] = 8'd154;
    assign expected_output[136] = 8'd128;
    assign expected_output[137] = 8'd154;
    assign expected_output[138] = 8'd228;
    assign expected_output[139] = 8'd58;
    assign expected_output[140] = 8'd126;
    assign expected_output[141] = 8'd127;
    assign expected_output[142] = 8'd127;
    assign expected_output[143] = 8'd127;
    assign expected_output[144] = 8'd126;
    assign expected_output[145] = 8'd127;
    assign expected_output[146] = 8'd127;
    assign expected_output[147] = 8'd127;
    assign expected_output[148] = 8'd127;
    assign expected_output[149] = 8'd58;
    assign expected_output[150] = 8'd224;
    assign expected_output[151] = 8'd150;
    assign expected_output[152] = 8'd128;
    assign expected_output[153] = 8'd170;
    assign expected_output[154] = 8'd4;
    assign expected_output[155] = 8'd90;
    assign expected_output[156] = 8'd126;
    assign expected_output[157] = 8'd90;
    assign expected_output[158] = 8'd4;
    assign expected_output[159] = 8'd170;
    assign expected_output[160] = 8'd128;
    assign expected_output[161] = 8'd150;
    assign expected_output[162] = 8'd224;
    assign expected_output[163] = 8'd58;
    assign expected_output[164] = 8'd124;
    assign expected_output[165] = 8'd127;
    assign expected_output[166] = 8'd127;
    assign expected_output[167] = 8'd127;
    assign expected_output[168] = 8'd127;
    assign expected_output[169] = 8'd120;
    assign expected_output[170] = 8'd116;
    assign expected_output[171] = 8'd120;
    assign expected_output[172] = 8'd124;
    assign expected_output[173] = 8'd127;
    assign expected_output[174] = 8'd127;
    assign expected_output[175] = 8'd127;
    assign expected_output[176] = 8'd127;
    assign expected_output[177] = 8'd58;
    assign expected_output[178] = 8'd224;
    assign expected_output[179] = 8'd150;
    assign expected_output[180] = 8'd128;
    assign expected_output[181] = 8'd170;
    assign expected_output[182] = 8'd4;
    assign expected_output[183] = 8'd90;
    assign expected_output[184] = 8'd127;
    assign expected_output[185] = 8'd90;
    assign expected_output[186] = 8'd0;
    assign expected_output[187] = 8'd166;
    assign expected_output[188] = 8'd130;
    assign expected_output[189] = 8'd166;
    assign expected_output[190] = 8'd252;
    assign expected_output[191] = 8'd86;
    assign expected_output[192] = 8'd126;
    assign expected_output[193] = 8'd106;
    assign expected_output[194] = 8'd36;
    assign expected_output[195] = 8'd202;
    assign expected_output[196] = 8'd132;
    assign expected_output[197] = 8'd128;
    assign expected_output[198] = 8'd128;
    assign expected_output[199] = 8'd128;
    assign expected_output[200] = 8'd128;
    assign expected_output[201] = 8'd202;
    assign expected_output[202] = 8'd36;
    assign expected_output[203] = 8'd106;
    assign expected_output[204] = 8'd127;
    assign expected_output[205] = 8'd86;
    assign expected_output[206] = 8'd0;
    assign expected_output[207] = 8'd170;
    assign expected_output[208] = 8'd130;
    assign expected_output[209] = 8'd150;
    assign expected_output[210] = 8'd220;
    assign expected_output[211] = 8'd54;
    assign expected_output[212] = 8'd126;
    assign expected_output[213] = 8'd127;
    assign expected_output[214] = 8'd127;
    assign expected_output[215] = 8'd127;
    assign expected_output[216] = 8'd127;
    assign expected_output[217] = 8'd70;
    assign expected_output[218] = 8'd252;
    assign expected_output[219] = 8'd182;
    assign expected_output[220] = 8'd130;
    assign expected_output[221] = 8'd128;
    assign expected_output[222] = 8'd128;
    assign expected_output[223] = 8'd128;
    assign expected_output[224] = 8'd130;
    assign expected_output[225] = 8'd136;
    assign expected_output[226] = 8'd136;
    assign expected_output[227] = 8'd132;
    assign expected_output[228] = 8'd132;
    assign expected_output[229] = 8'd132;
    assign expected_output[230] = 8'd132;
    assign expected_output[231] = 8'd132;
    assign expected_output[232] = 8'd130;
    assign expected_output[233] = 8'd132;
    assign expected_output[234] = 8'd136;
    assign expected_output[235] = 8'd136;
    assign expected_output[236] = 8'd132;
    assign expected_output[237] = 8'd128;
    assign expected_output[238] = 8'd128;
    assign expected_output[239] = 8'd128;
    assign expected_output[240] = 8'd130;
    assign expected_output[241] = 8'd198;
    assign expected_output[242] = 8'd28;
    assign expected_output[243] = 8'd102;
    assign expected_output[244] = 8'd127;
    assign expected_output[245] = 8'd102;
    assign expected_output[246] = 8'd32;
    assign expected_output[247] = 8'd202;
    assign expected_output[248] = 8'd130;
    assign expected_output[249] = 8'd128;
    assign expected_output[250] = 8'd128;
    assign expected_output[251] = 8'd128;
    assign expected_output[252] = 8'd128;
    assign expected_output[253] = 8'd186;
    assign expected_output[254] = 8'd0;
    assign expected_output[255] = 8'd70;
    assign expected_output[256] = 8'd126;
    assign expected_output[257] = 8'd127;
    assign expected_output[258] = 8'd127;
    assign expected_output[259] = 8'd127;
    assign expected_output[260] = 8'd127;
    assign expected_output[261] = 8'd54;
    assign expected_output[262] = 8'd224;
    assign expected_output[263] = 8'd154;
    assign expected_output[264] = 8'd128;
    assign expected_output[265] = 8'd154;
    assign expected_output[266] = 8'd224;
    assign expected_output[267] = 8'd54;
    assign expected_output[268] = 8'd124;
    assign expected_output[269] = 8'd127;
    assign expected_output[270] = 8'd127;
    assign expected_output[271] = 8'd127;
    assign expected_output[272] = 8'd127;
    assign expected_output[273] = 8'd54;
    assign expected_output[274] = 8'd224;
    assign expected_output[275] = 8'd154;
    assign expected_output[276] = 8'd128;
    assign expected_output[277] = 8'd154;
    assign expected_output[278] = 8'd224;
    assign expected_output[279] = 8'd54;
    assign expected_output[280] = 8'd124;
    assign expected_output[281] = 8'd127;
    assign expected_output[282] = 8'd127;
    assign expected_output[283] = 8'd127;
    assign expected_output[284] = 8'd127;
    assign expected_output[285] = 8'd54;
    assign expected_output[286] = 8'd220;
    assign expected_output[287] = 8'd150;
    assign expected_output[288] = 8'd128;
    assign expected_output[289] = 8'd170;
    assign expected_output[290] = 8'd0;
    assign expected_output[291] = 8'd86;
    assign expected_output[292] = 8'd126;
    assign expected_output[293] = 8'd106;
    assign expected_output[294] = 8'd36;
    assign expected_output[295] = 8'd202;
    assign expected_output[296] = 8'd132;
    assign expected_output[297] = 8'd128;
    assign expected_output[298] = 8'd128;
    assign expected_output[299] = 8'd128;
    assign expected_output[300] = 8'd128;
    assign expected_output[301] = 8'd202;
    assign expected_output[302] = 8'd32;
    assign expected_output[303] = 8'd102;
    assign expected_output[304] = 8'd127;
    assign expected_output[305] = 8'd102;
    assign expected_output[306] = 8'd28;
    assign expected_output[307] = 8'd198;
    assign expected_output[308] = 8'd132;
    assign expected_output[309] = 8'd128;
    assign expected_output[310] = 8'd128;
    assign expected_output[311] = 8'd128;
    assign expected_output[312] = 8'd130;
    assign expected_output[313] = 8'd136;
    assign expected_output[314] = 8'd136;
    assign expected_output[315] = 8'd132;
    assign expected_output[316] = 8'd132;
    assign expected_output[317] = 8'd132;
    assign expected_output[318] = 8'd132;
    assign expected_output[319] = 8'd132;
    assign expected_output[320] = 8'd130;
    assign expected_output[321] = 8'd132;
    assign expected_output[322] = 8'd136;
    assign expected_output[323] = 8'd136;
    assign expected_output[324] = 8'd130;
    assign expected_output[325] = 8'd128;
    assign expected_output[326] = 8'd128;
    assign expected_output[327] = 8'd128;
    assign expected_output[328] = 8'd130;
    assign expected_output[329] = 8'd182;
    assign expected_output[330] = 8'd252;
    assign expected_output[331] = 8'd70;
    assign expected_output[332] = 8'd126;
    assign expected_output[333] = 8'd127;
    assign expected_output[334] = 8'd127;
    assign expected_output[335] = 8'd127;
    assign expected_output[336] = 8'd127;
    assign expected_output[337] = 8'd54;
    assign expected_output[338] = 8'd224;
    assign expected_output[339] = 8'd154;
    assign expected_output[340] = 8'd128;
    assign expected_output[341] = 8'd154;
    assign expected_output[342] = 8'd224;
    assign expected_output[343] = 8'd54;
    assign expected_output[344] = 8'd126;
    assign expected_output[345] = 8'd127;
    assign expected_output[346] = 8'd127;
    assign expected_output[347] = 8'd127;
    assign expected_output[348] = 8'd127;
    assign expected_output[349] = 8'd70;
    assign expected_output[350] = 8'd0;
    assign expected_output[351] = 8'd186;
    assign expected_output[352] = 8'd130;
    assign expected_output[353] = 8'd128;
    assign expected_output[354] = 8'd128;
    assign expected_output[355] = 8'd128;
    assign expected_output[356] = 8'd128;
    assign expected_output[357] = 8'd202;
    assign expected_output[358] = 8'd36;
    assign expected_output[359] = 8'd106;
    assign expected_output[360] = 8'd127;
    assign expected_output[361] = 8'd86;
    assign expected_output[362] = 8'd252;
    assign expected_output[363] = 8'd166;
    assign expected_output[364] = 8'd128;
    assign expected_output[365] = 8'd166;
    assign expected_output[366] = 8'd0;
    assign expected_output[367] = 8'd90;
    assign expected_output[368] = 8'd126;
    assign expected_output[369] = 8'd90;
    assign expected_output[370] = 8'd4;
    assign expected_output[371] = 8'd170;
    assign expected_output[372] = 8'd130;
    assign expected_output[373] = 8'd150;
    assign expected_output[374] = 8'd220;
    assign expected_output[375] = 8'd54;
    assign expected_output[376] = 8'd126;
    assign expected_output[377] = 8'd127;
    assign expected_output[378] = 8'd127;
    assign expected_output[379] = 8'd127;
    assign expected_output[380] = 8'd127;
    assign expected_output[381] = 8'd70;
    assign expected_output[382] = 8'd0;
    assign expected_output[383] = 8'd186;
    assign expected_output[384] = 8'd128;
    assign expected_output[385] = 8'd128;
    assign expected_output[386] = 8'd128;
    assign expected_output[387] = 8'd128;
    assign expected_output[388] = 8'd128;
    assign expected_output[389] = 8'd186;
    assign expected_output[390] = 8'd0;
    assign expected_output[391] = 8'd70;
    assign expected_output[392] = 8'd127;
    assign expected_output[393] = 8'd127;
    assign expected_output[394] = 8'd127;
    assign expected_output[395] = 8'd127;
    assign expected_output[396] = 8'd127;
    assign expected_output[397] = 8'd70;
    assign expected_output[398] = 8'd0;
    assign expected_output[399] = 8'd186;
    assign expected_output[400] = 8'd128;
    assign expected_output[401] = 8'd128;
    assign expected_output[402] = 8'd128;
    assign expected_output[403] = 8'd128;
    assign expected_output[404] = 8'd128;
    assign expected_output[405] = 8'd186;
    assign expected_output[406] = 8'd4;
    assign expected_output[407] = 8'd74;
    assign expected_output[408] = 8'd126;
    assign expected_output[409] = 8'd127;
    assign expected_output[410] = 8'd127;
    assign expected_output[411] = 8'd127;
    assign expected_output[412] = 8'd126;
    assign expected_output[413] = 8'd120;
    assign expected_output[414] = 8'd120;
    assign expected_output[415] = 8'd124;
    assign expected_output[416] = 8'd124;
    assign expected_output[417] = 8'd124;
    assign expected_output[418] = 8'd124;
    assign expected_output[419] = 8'd124;
    assign expected_output[420] = 8'd124;
    assign expected_output[421] = 8'd124;
    assign expected_output[422] = 8'd124;
    assign expected_output[423] = 8'd124;
    assign expected_output[424] = 8'd126;
    assign expected_output[425] = 8'd124;
    assign expected_output[426] = 8'd120;
    assign expected_output[427] = 8'd120;
    assign expected_output[428] = 8'd126;
    assign expected_output[429] = 8'd127;
    assign expected_output[430] = 8'd127;
    assign expected_output[431] = 8'd127;
    assign expected_output[432] = 8'd126;
    assign expected_output[433] = 8'd74;
    assign expected_output[434] = 8'd4;
    assign expected_output[435] = 8'd186;
    assign expected_output[436] = 8'd128;
    assign expected_output[437] = 8'd128;
    assign expected_output[438] = 8'd128;
    assign expected_output[439] = 8'd128;
    assign expected_output[440] = 8'd128;
    assign expected_output[441] = 8'd186;
    assign expected_output[442] = 8'd4;
    assign expected_output[443] = 8'd74;
    assign expected_output[444] = 8'd127;
    assign expected_output[445] = 8'd127;
    assign expected_output[446] = 8'd127;
    assign expected_output[447] = 8'd127;
    assign expected_output[448] = 8'd127;
    assign expected_output[449] = 8'd127;
    assign expected_output[450] = 8'd127;
    assign expected_output[451] = 8'd127;
    assign expected_output[452] = 8'd126;
    assign expected_output[453] = 8'd74;
    assign expected_output[454] = 8'd4;
    assign expected_output[455] = 8'd186;
    assign expected_output[456] = 8'd128;
    assign expected_output[457] = 8'd128;
    assign expected_output[458] = 8'd128;
    assign expected_output[459] = 8'd128;
    assign expected_output[460] = 8'd128;
    assign expected_output[461] = 8'd186;
    assign expected_output[462] = 8'd0;
    assign expected_output[463] = 8'd70;
    assign expected_output[464] = 8'd126;
    assign expected_output[465] = 8'd127;
    assign expected_output[466] = 8'd127;
    assign expected_output[467] = 8'd127;
    assign expected_output[468] = 8'd127;
    assign expected_output[469] = 8'd54;
    assign expected_output[470] = 8'd220;
    assign expected_output[471] = 8'd150;
    assign expected_output[472] = 8'd128;
    assign expected_output[473] = 8'd170;
    assign expected_output[474] = 8'd4;
    assign expected_output[475] = 8'd90;
    assign expected_output[476] = 8'd126;
    assign expected_output[477] = 8'd90;
    assign expected_output[478] = 8'd4;
    assign expected_output[479] = 8'd170;
    assign expected_output[480] = 8'd128;
    assign expected_output[481] = 8'd150;
    assign expected_output[482] = 8'd224;
    assign expected_output[483] = 8'd58;
    assign expected_output[484] = 8'd126;
    assign expected_output[485] = 8'd127;
    assign expected_output[486] = 8'd127;
    assign expected_output[487] = 8'd127;
    assign expected_output[488] = 8'd127;
    assign expected_output[489] = 8'd127;
    assign expected_output[490] = 8'd127;
    assign expected_output[491] = 8'd127;
    assign expected_output[492] = 8'd126;
    assign expected_output[493] = 8'd74;
    assign expected_output[494] = 8'd4;
    assign expected_output[495] = 8'd186;
    assign expected_output[496] = 8'd130;
    assign expected_output[497] = 8'd128;
    assign expected_output[498] = 8'd128;
    assign expected_output[499] = 8'd128;
    assign expected_output[500] = 8'd128;
    assign expected_output[501] = 8'd202;
    assign expected_output[502] = 8'd36;
    assign expected_output[503] = 8'd106;
    assign expected_output[504] = 8'd127;
    assign expected_output[505] = 8'd86;
    assign expected_output[506] = 8'd0;
    assign expected_output[507] = 8'd170;
    assign expected_output[508] = 8'd130;
    assign expected_output[509] = 8'd150;
    assign expected_output[510] = 8'd220;
    assign expected_output[511] = 8'd54;
    assign expected_output[512] = 8'd124;
    assign expected_output[513] = 8'd127;
    assign expected_output[514] = 8'd127;
    assign expected_output[515] = 8'd127;
    assign expected_output[516] = 8'd127;
    assign expected_output[517] = 8'd54;
    assign expected_output[518] = 8'd220;
    assign expected_output[519] = 8'd150;
    assign expected_output[520] = 8'd128;
    assign expected_output[521] = 8'd170;
    assign expected_output[522] = 8'd0;
    assign expected_output[523] = 8'd86;
    assign expected_output[524] = 8'd127;
    assign expected_output[525] = 8'd106;
    assign expected_output[526] = 8'd32;
    assign expected_output[527] = 8'd198;
    assign expected_output[528] = 8'd132;
    assign expected_output[529] = 8'd128;
    assign expected_output[530] = 8'd128;
    assign expected_output[531] = 8'd128;
    assign expected_output[532] = 8'd130;
    assign expected_output[533] = 8'd136;
    assign expected_output[534] = 8'd136;
    assign expected_output[535] = 8'd132;
    assign expected_output[536] = 8'd132;
    assign expected_output[537] = 8'd132;
    assign expected_output[538] = 8'd132;
    assign expected_output[539] = 8'd132;
    assign expected_output[540] = 8'd132;
    assign expected_output[541] = 8'd132;
    assign expected_output[542] = 8'd132;
    assign expected_output[543] = 8'd132;
    assign expected_output[544] = 8'd130;
    assign expected_output[545] = 8'd132;
    assign expected_output[546] = 8'd136;
    assign expected_output[547] = 8'd136;
    assign expected_output[548] = 8'd132;
    assign expected_output[549] = 8'd128;
    assign expected_output[550] = 8'd128;
    assign expected_output[551] = 8'd128;
    assign expected_output[552] = 8'd128;
    assign expected_output[553] = 8'd198;
    assign expected_output[554] = 8'd32;
    assign expected_output[555] = 8'd106;
    assign expected_output[556] = 8'd127;
    assign expected_output[557] = 8'd86;
    assign expected_output[558] = 8'd0;
    assign expected_output[559] = 8'd170;
    assign expected_output[560] = 8'd128;
    assign expected_output[561] = 8'd150;
    assign expected_output[562] = 8'd224;
    assign expected_output[563] = 8'd58;
    assign expected_output[564] = 8'd126;
    assign expected_output[565] = 8'd127;
    assign expected_output[566] = 8'd127;
    assign expected_output[567] = 8'd127;
    assign expected_output[568] = 8'd126;
    assign expected_output[569] = 8'd127;
    assign expected_output[570] = 8'd127;
    assign expected_output[571] = 8'd127;
    assign expected_output[572] = 8'd127;
    assign expected_output[573] = 8'd58;
    assign expected_output[574] = 8'd224;
    assign expected_output[575] = 8'd150;
    assign expected_output[576] = 8'd128;
    assign expected_output[577] = 8'd170;
    assign expected_output[578] = 8'd0;
    assign expected_output[579] = 8'd86;
    assign expected_output[580] = 8'd126;
    assign expected_output[581] = 8'd106;
    assign expected_output[582] = 8'd36;
    assign expected_output[583] = 8'd202;
    assign expected_output[584] = 8'd130;
    assign expected_output[585] = 8'd128;
    assign expected_output[586] = 8'd128;
    assign expected_output[587] = 8'd128;
    assign expected_output[588] = 8'd128;
    assign expected_output[589] = 8'd186;
    assign expected_output[590] = 8'd4;
    assign expected_output[591] = 8'd74;
    assign expected_output[592] = 8'd127;
    assign expected_output[593] = 8'd127;
    assign expected_output[594] = 8'd127;
    assign expected_output[595] = 8'd127;
    assign expected_output[596] = 8'd127;
    assign expected_output[597] = 8'd127;
    assign expected_output[598] = 8'd127;
    assign expected_output[599] = 8'd127;
    assign expected_output[600] = 8'd127;
    assign expected_output[601] = 8'd74;
    assign expected_output[602] = 8'd0;
    assign expected_output[603] = 8'd182;
    assign expected_output[604] = 8'd128;
    assign expected_output[605] = 8'd128;
    assign expected_output[606] = 8'd128;
    assign expected_output[607] = 8'd128;
    assign expected_output[608] = 8'd130;
    assign expected_output[609] = 8'd128;
    assign expected_output[610] = 8'd128;
    assign expected_output[611] = 8'd128;
    assign expected_output[612] = 8'd128;
    assign expected_output[613] = 8'd198;
    assign expected_output[614] = 8'd32;
    assign expected_output[615] = 8'd106;
    assign expected_output[616] = 8'd127;
    assign expected_output[617] = 8'd86;
    assign expected_output[618] = 8'd252;
    assign expected_output[619] = 8'd166;
    assign expected_output[620] = 8'd130;
    assign expected_output[621] = 8'd166;
    assign expected_output[622] = 8'd252;
    assign expected_output[623] = 8'd86;
    assign expected_output[624] = 8'd126;
    assign expected_output[625] = 8'd106;
    assign expected_output[626] = 8'd36;
    assign expected_output[627] = 8'd202;
    assign expected_output[628] = 8'd130;
    assign expected_output[629] = 8'd128;
    assign expected_output[630] = 8'd128;
    assign expected_output[631] = 8'd128;
    assign expected_output[632] = 8'd128;
    assign expected_output[633] = 8'd186;
    assign expected_output[634] = 8'd0;
    assign expected_output[635] = 8'd70;
    assign expected_output[636] = 8'd126;
    assign expected_output[637] = 8'd127;
    assign expected_output[638] = 8'd127;
    assign expected_output[639] = 8'd127;
    assign expected_output[640] = 8'd127;
    assign expected_output[641] = 8'd54;
    assign expected_output[642] = 8'd220;
    assign expected_output[643] = 8'd150;
    assign expected_output[644] = 8'd128;
    assign expected_output[645] = 8'd170;
    assign expected_output[646] = 8'd0;
    assign expected_output[647] = 8'd86;
    assign expected_output[648] = 8'd126;
    assign expected_output[649] = 8'd106;
    assign expected_output[650] = 8'd36;
    assign expected_output[651] = 8'd202;
    assign expected_output[652] = 8'd130;
    assign expected_output[653] = 8'd128;
    assign expected_output[654] = 8'd128;
    assign expected_output[655] = 8'd128;
    assign expected_output[656] = 8'd128;
    assign expected_output[657] = 8'd186;
    assign expected_output[658] = 8'd0;
    assign expected_output[659] = 8'd70;
    assign expected_output[660] = 8'd127;
    assign expected_output[661] = 8'd127;
    assign expected_output[662] = 8'd127;
    assign expected_output[663] = 8'd127;
    assign expected_output[664] = 8'd127;
    assign expected_output[665] = 8'd70;
    assign expected_output[666] = 8'd252;
    assign expected_output[667] = 8'd182;
    assign expected_output[668] = 8'd130;
    assign expected_output[669] = 8'd128;
    assign expected_output[670] = 8'd128;
    assign expected_output[671] = 8'd128;
    assign expected_output[672] = 8'd128;
    assign expected_output[673] = 8'd136;
    assign expected_output[674] = 8'd140;
    assign expected_output[675] = 8'd136;
    assign expected_output[676] = 8'd130;
    assign expected_output[677] = 8'd128;
    assign expected_output[678] = 8'd128;
    assign expected_output[679] = 8'd128;
    assign expected_output[680] = 8'd128;
    assign expected_output[681] = 8'd182;
    assign expected_output[682] = 8'd0;
    assign expected_output[683] = 8'd74;
    assign expected_output[684] = 8'd127;
    assign expected_output[685] = 8'd127;
    assign expected_output[686] = 8'd127;
    assign expected_output[687] = 8'd127;
    assign expected_output[688] = 8'd127;
    assign expected_output[689] = 8'd127;
    assign expected_output[690] = 8'd127;
    assign expected_output[691] = 8'd127;
    assign expected_output[692] = 8'd127;
    assign expected_output[693] = 8'd74;
    assign expected_output[694] = 8'd0;
    assign expected_output[695] = 8'd182;
    assign expected_output[696] = 8'd130;
    assign expected_output[697] = 8'd128;
    assign expected_output[698] = 8'd128;
    assign expected_output[699] = 8'd128;
    assign expected_output[700] = 8'd130;
    assign expected_output[701] = 8'd136;
    assign expected_output[702] = 8'd136;
    assign expected_output[703] = 8'd132;
    assign expected_output[704] = 8'd130;
    assign expected_output[705] = 8'd132;
    assign expected_output[706] = 8'd136;
    assign expected_output[707] = 8'd136;
    assign expected_output[708] = 8'd132;
    assign expected_output[709] = 8'd128;
    assign expected_output[710] = 8'd128;
    assign expected_output[711] = 8'd128;
    assign expected_output[712] = 8'd130;
    assign expected_output[713] = 8'd198;
    assign expected_output[714] = 8'd28;
    assign expected_output[715] = 8'd102;
    assign expected_output[716] = 8'd127;
    assign expected_output[717] = 8'd102;
    assign expected_output[718] = 8'd28;
    assign expected_output[719] = 8'd198;
    assign expected_output[720] = 8'd130;
    assign expected_output[721] = 8'd128;
    assign expected_output[722] = 8'd128;
    assign expected_output[723] = 8'd128;
    assign expected_output[724] = 8'd130;
    assign expected_output[725] = 8'd128;
    assign expected_output[726] = 8'd128;
    assign expected_output[727] = 8'd128;
    assign expected_output[728] = 8'd128;
    assign expected_output[729] = 8'd198;
    assign expected_output[730] = 8'd32;
    assign expected_output[731] = 8'd106;
    assign expected_output[732] = 8'd127;
    assign expected_output[733] = 8'd86;
    assign expected_output[734] = 8'd0;
    assign expected_output[735] = 8'd170;
    assign expected_output[736] = 8'd128;
    assign expected_output[737] = 8'd150;
    assign expected_output[738] = 8'd224;
    assign expected_output[739] = 8'd58;
    assign expected_output[740] = 8'd124;
    assign expected_output[741] = 8'd127;
    assign expected_output[742] = 8'd127;
    assign expected_output[743] = 8'd127;
    assign expected_output[744] = 8'd126;
    assign expected_output[745] = 8'd120;
    assign expected_output[746] = 8'd120;
    assign expected_output[747] = 8'd124;
    assign expected_output[748] = 8'd126;
    assign expected_output[749] = 8'd124;
    assign expected_output[750] = 8'd120;
    assign expected_output[751] = 8'd120;
    assign expected_output[752] = 8'd126;
    assign expected_output[753] = 8'd127;
    assign expected_output[754] = 8'd127;
    assign expected_output[755] = 8'd127;
    assign expected_output[756] = 8'd126;
    assign expected_output[757] = 8'd74;
    assign expected_output[758] = 8'd4;
    assign expected_output[759] = 8'd186;
    assign expected_output[760] = 8'd130;
    assign expected_output[761] = 8'd128;
    assign expected_output[762] = 8'd128;
    assign expected_output[763] = 8'd128;
    assign expected_output[764] = 8'd128;
    assign expected_output[765] = 8'd202;
    assign expected_output[766] = 8'd36;
    assign expected_output[767] = 8'd106;
    assign expected_output[768] = 8'd127;
    assign expected_output[769] = 8'd86;
    assign expected_output[770] = 8'd252;
    assign expected_output[771] = 8'd166;
    assign expected_output[772] = 8'd130;
    assign expected_output[773] = 8'd166;
    assign expected_output[774] = 8'd252;
    assign expected_output[775] = 8'd86;
    assign expected_output[776] = 8'd126;
    assign expected_output[777] = 8'd106;
    assign expected_output[778] = 8'd36;
    assign expected_output[779] = 8'd202;
    assign expected_output[780] = 8'd132;
    assign expected_output[781] = 8'd128;
    assign expected_output[782] = 8'd128;
    assign expected_output[783] = 8'd128;
    assign expected_output[784] = 8'd128;
    assign expected_output[785] = 8'd202;
    assign expected_output[786] = 8'd32;
    assign expected_output[787] = 8'd102;
    assign expected_output[788] = 8'd127;
    assign expected_output[789] = 8'd102;
    assign expected_output[790] = 8'd32;
    assign expected_output[791] = 8'd202;
    assign expected_output[792] = 8'd132;
    assign expected_output[793] = 8'd128;
    assign expected_output[794] = 8'd128;
    assign expected_output[795] = 8'd128;
    assign expected_output[796] = 8'd128;
    assign expected_output[797] = 8'd202;
    assign expected_output[798] = 8'd32;
    assign expected_output[799] = 8'd102;
endmodule